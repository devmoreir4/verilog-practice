module CodTeclado (tecla, cod_gray);
	
	input [3:0] tecla;
	output [3:0] cod_gray;
	
endmodule 